/*-----------------------------------------------------------------
taylor.templeton@gmail.com
May 2023

Verification Practice Project
Verify each block -> Verify CPU
-----------------------------------------------------------------*/
package testbench_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "sequence_items.sv"
`include "sequencer.sv"
`include "sequence.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "scoreboard.sv"
`include "functional_coverage.sv"
`include "environment.sv"
`include "test.sv"

endpackage : testbench_pkg